// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module adder(
    input  A,
    input  B,
    input Clk,
    input En,
    output [3:0] Sum,
    output Overflow
    );
    
endmodule